module main

struct AuthRequestDto{
	username string [required]
	password string [required]
}